module	
	

endmodule
